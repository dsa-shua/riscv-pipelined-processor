`timescale 1ns / 1ps
module AND_GATE(
    input A,B,
    output wire C
    );
    
    assign C = A & B;
endmodule
