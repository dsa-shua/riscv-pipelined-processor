module controller(
    output wire [31:0] r0,
    output wire [31:0] r1,
    output wire [31:0] r2,
    output wire [31:0] r3,
    output wire [31:0] r4,
    output wire [31:0] r5,
    output wire [31:0] r6,
    output wire [31:0] r7
    
);
    assign r0 = 32'd15;
    assign r1 = 32'd7;
    assign r2 = 32'd18;
    assign r3 = 32'd55;
    assign r4 = 32'd42;
    assign r5 = 32'd17;
    assign r6 = 32'd5;
    assign r7 = 32'd81;
   
    
endmodule